0
0 6 0 9 0r 38 47 43 h 37 T 25 T 30 B
0 2 0 0 0r 56 48 64 h 32 H 44 B
11 0 0 0 0r 24 50 33 41 h 16 H 40 B
0 0 3 0 0r 27 32 h 20 H 27 H
BRICK 3ENERGY 10HEAT 5ENERGY 4PARK 7HEAT 10GLASS 11BRICK 3HEAT 8BRICK 2BRICK 6ENERGY 8WIFI 12ENERGY 5WIFI 11GLASS 4WIFI 6GLASS 9GLASS 9
7
